// file: ForwardUnit.v
// author: @mobs_11

`timescale 1ns/1ns

module ForwardUnit;

endmodule